----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:16:25 12/01/2016 
-- Design Name: 
-- Module Name:    mux2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2 is
    Port ( 
			  rt 		: IN  	STD_LOGIC_VECTOR (31 downto 0);
           imm 	: IN  	STD_LOGIC_VECTOR (31 downto 0);
			  sel 	: IN 		STD_LOGIC;
           output : OUT  	STD_LOGIC_VECTOR (31 downto 0)
			 );
end mux2;

architecture Behavioral of mux2 is

begin

WITH sel SELECT 
	output <= rt WHEN '0',
				 imm WHEN '1';

end Behavioral;

