----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:23:23 11/27/2016 
-- Design Name: 
-- Module Name:    instr_mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity instr_mem is
	PORT 
	(		
		clr			: IN STD_LOGIC;
		read_addr	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		instr		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	 );
end instr_mem;

architecture Behavioral of instr_mem is
	
	constant DATA_BITS : Integer := 32;			-- no of bits per word
	constant DEPTH     : Integer := 256;		-- no of lines TODO change depth to 2 power 32
--	constant FILENAME  : String(1 to 19) := "inputfilename.hex";
	
	
	subtype word_t  is std_logic_vector(DATA_BITS - 1 downto 0);
	type    ram_t   is array(0 to DEPTH - 1) of word_t;
--	signal ram    : ram_t    := ReadAssemblyFile(FILENAME);
	signal ram    : ram_t := 	(X"00000000",	
"00000100000000110000000000000100",
"00000100000000010000000000000001",
"00001000011000110000000000000001",
"00011100011000100000000000000000",
"00100000011000100000000000001010",
"00101100000000111111111111111100",
"00011100000000100000000000001000",
"00100000000000100000000000001110",
"00011100000001000000000000001001",
"00000100000001110000000000011011",
"00000000100000100001000000010000",
"00100000001000100000000000001110",
"00000100001000010000000000000001",
"00101100111000011111111111111100",
"00000100000000010000000000000000",
"00000100001000100000000000000000",
"00000100001000110000000000000000",
"00000100001001000000000000000000",
"00000100001001010000000000000000",
"00000100000010000000000000000100",
"00000100000010010000000001001110",
"00000100000100000000000000011010",
"00011100001001100000000000001110",
"00000000100000110001100000010000",
"00000000110000110001100000010000",
"00000100000010110000000000000011",
"00100000000000110000000000110000",
"00100000000010110000000000110001",
"00000101011010111111111111111101",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00010101011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00011001111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00100000001010110000000000001110",
"00000001011000000001100000010000",
"00011100010001100000000000001010",
"00000100100001000000000000000000",
"00000000100000111010000000010000",
"00000000110101000010000000010000",
"00100000000001000000000000110000",
"00100000000101000000000000110001",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00010101011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00011001111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00100000010010110000000000001010",
"00000001011000000010000000010000",
"00000100001000010000000000000001",
"00000100010000100000000000000001",
"00101110000000010000000000000001",
"00000100000000010000000000000000",
"00101101000000100000000000000001",
"00000100000000100000000000000000",
"00000100101001010000000000000001",
"00101101001001011111111111001011",
"00000100000000010000000000000000",
"00011100001000100000000000001110",
"00011100001000110000000000101011",
"00000000011000100001100000010000",
"00000100001000010000000000000001",
"00011100001001000000000000001110",
"00011100001001010000000000101011",
"00000000101001000010100000010000",
"00000100000101000000000000001101",
"00000100001010000000000000000000",
"00000000101000110011000000010010",
"00000000101000110011100000010100",
"00000000111001100011100000010100",
"00100000000001110000000000110000",
"00100000000001010000000000110001",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00010101011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00011001111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00000001000010000100000000010000",
"00011101000010010000000000001110",
"00000001001010110001100000010000",
"00000100011000110000000000000000",
"00000000101000110011000000010010",
"00000000101000110011100000010100",
"00000000111001100011100000010100",
"00100000000001110000000000110000",
"00100000000000110000000000110001",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00010101011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00011001111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00000101000010000000000000000001",
"00011101000010010000000000001110",
"00000001001010110010100000010000",
"00000100101001010000000000000000",
"00000100001000010000000000000001",
"00101110100000011111111111010010",
"00000100000000010000000000000000",
"00100000001000110000000000101101",
"00000100011000110000000000000000",
"00000100001000010000000000000001",
"00100000001001010000000000101101",
"00000100101001010000000000000000",
"00000100000000010000000000000000",
"00011100001000110000000000101101",
"00000100001000010000000000000001",
"00011100001001010000000000101101",
"00000100000100000000000000000001",
"00000100000000010000000000001100",
"00000100001000100000000000000000",
"00000000001000010000100000010000",
"00000100001000010000000000000001",
"00011100001001100000000000001110",
"00000000110001010010100000010001",
"00100000000001010000000000110000",
"00100000000000110000000000110001",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00011001011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00010101111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00000000011010110100000000010010",
"00000000011010110011100000010100",
"00000000111010000010100000010100",
"00001000001000010000000000000001",
"00011100001001100000000000001110",
"00000000110000110001100000010001",
"00100000000000110000000000110000",
"00100000000001010000000000110001",
"00011100000010100000000000101111",
"00011100000010110000000000110000",
"00011100000011000000000000110001",
"00000001010011000110100000010010",
"00101000000011010000000000001001",
"00001001101011100000000000100000",
"00011100000011110000000000110000",
"00011001011010110000000000000001",
"00001001101011010000000000000001",
"00101100000011011111111111111101",
"00010101111011110000000000000001",
"00000101110011100000000000000001",
"00101100000011101111111111111101",
"00000001111010110101100000010011",
"00000000101010110100000000010010",
"00000000101010110011100000010100",
"00000000111010000001100000010100",
"00001000001000010000000000000001",
"00101110000000011111111111010010",
"00011100001001100000000000001110",
"00000000110001010010100000010001",
"00001000001000010000000000000001",
"00011100001001100000000000001110",
"00000000110000110001100000010001",
"00100000000000110000000000101011",
"00000100011000110000000000000000",
"00100000000001010000000000101100",
"00000100101001010000000000000000",			
"11111100000000000000000000000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00000000",X"00000000",X"00000000",X"00000000");
	
	
	-- Read a *.hex file
	-- TODO hard code the values into instruction memory
--	impure function ReadBinaryFile(FileName : STRING) return ram_t is
--		file FileHandle       : TEXT open READ_MODE is FileName;
--		variable CurrentLine  : LINE;
--		variable TempWord     : STD_LOGIC_VECTOR((div_ceil(word_t'length, 4) * 4) - 1 downto 0);
--		variable Result       : ram_t    := (others => (others => '0'));
--
--		begin
--		for i in 0 to DEPTH - 1 loop
--		 exit when endfile(FileHandle);
--
--		 readline(FileHandle, CurrentLine);
--		 hread(CurrentLine, TempWord);
--		 Result(i)    := resize(TempWord, word_t'length);
--		end loop;
--
--		return Result;
--	end function;
	
	
begin


	PROCESS(clr)
	BEGIN
		IF (clr = '1') THEN
		null;
--ram(1) <= "00000100000000110000000000000100";
--ram(2) <= "00000100000000010000000000000001";
--ram(3) <= "00001000011000110000000000000001";
--ram(4) <= "00011100011000100000000000000000";
--ram(5) <= "00100000011000100000000000001010";
--ram(6) <= "00101100000000111111111111111100";
--ram(7) <= "00011100000000100000000000001000";
--ram(8) <= "00100000000000100000000000001110";
--ram(9) <= "00011100000001000000000000001001";
--ram(10) <= "00000100000001110000000000011011";
--ram(11) <= "00000000100000100001000000010000";
--ram(12) <= "00100000001000100000000000001110";
--ram(13) <= "00000100001000010000000000000001";
--ram(14) <= "00101100111000011111111111111100";
--ram(15) <= "00000100000000010000000000000000";
--ram(16) <= "00000100001000100000000000000000";
--ram(17) <= "00000100001000110000000000000000";
--ram(18) <= "00000100001001000000000000000000";
--ram(19) <= "00000100001001010000000000000000";
--ram(20) <= "00000100000010000000000000000100";
--ram(21) <= "00000100000010010000000001001110";
--ram(22) <= "00000100000100000000000000011010";
--ram(23) <= "00011100001001100000000000001110";
--ram(24) <= "00000000100000110001100000010000";
--ram(25) <= "00000000110000110001100000010000";
--ram(26) <= "00000100000010110000000000000011";
--ram(27) <= "00100000000000110000000000110000";
--ram(28) <= "00100000000010110000000000110001";
--ram(29) <= "00000101011010111111111111111101";
--ram(30) <= "00011100000010100000000000101111";
--ram(31) <= "00011100000010110000000000110000";
--ram(32) <= "00011100000011000000000000110001";
--ram(33) <= "00000001010011000110100000010010";
--ram(34) <= "00101000000011010000000000001001";
--ram(35) <= "00001001101011100000000000100000";
--ram(36) <= "00011100000011110000000000110000";
--ram(37) <= "00010101011010110000000000000001";
--ram(38) <= "00001001101011010000000000000001";
--ram(39) <= "00101100000011011111111111111101";
--ram(40) <= "00011001111011110000000000000001";
--ram(41) <= "00000101110011100000000000000001";
--ram(42) <= "00101100000011101111111111111101";
--ram(43) <= "00000001111010110101100000010011";
--ram(44) <= "00100000001010110000000000001110";
--ram(45) <= "00000001011000000001100000010000";
--ram(46) <= "00011100010001100000000000001010";
--ram(47) <= "00000100100001000000000000000000";
--ram(48) <= "00000000100000111010000000010000";
--ram(49) <= "00000000110101000010000000010000";
--ram(50) <= "00100000000001000000000000110000";
--ram(51) <= "00100000000101000000000000110001";
--ram(52) <= "00011100000010100000000000101111";
--ram(53) <= "00011100000010110000000000110000";
--ram(54) <= "00011100000011000000000000110001";
--ram(55) <= "00000001010011000110100000010010";
--ram(56) <= "00101000000011010000000000001001";
--ram(57) <= "00001001101011100000000000100000";
--ram(58) <= "00011100000011110000000000110000";
--ram(59) <= "00010101011010110000000000000001";
--ram(60) <= "00001001101011010000000000000001";
--ram(61) <= "00101100000011011111111111111101";
--ram(62) <= "00011001111011110000000000000001";
--ram(63) <= "00000101110011100000000000000001";
--ram(64) <= "00101100000011101111111111111101";
--ram(65) <= "00000001111010110101100000010011";
--ram(66) <= "00100000010010110000000000001010";
--ram(67) <= "00000001011000000010000000010000";
--ram(68) <= "00000100001000010000000000000001";
--ram(69) <= "00000100010000100000000000000001";
--ram(70) <= "00101110000000010000000000000001";
--ram(71) <= "00000100000000010000000000000000";
--ram(72) <= "00101101000000100000000000000001";
--ram(73) <= "00000100000000100000000000000000";
--ram(74) <= "00000100101001010000000000000001";
--ram(75) <= "00101101001001011111111111001011";
--ram(76) <= "00000100000000010000000000000000";
--ram(77) <= "00011100001000100000000000001110";
--ram(78) <= "00011100001000110000000000101011";
--ram(79) <= "00000000011000100001100000010000";
--ram(80) <= "00000100001000010000000000000001";
--ram(81) <= "00011100001001000000000000001110";
--ram(82) <= "00011100001001010000000000101011";
--ram(83) <= "00000000101001000010100000010000";
--ram(84) <= "00000100000101000000000000001101";
--ram(85) <= "00000100001010000000000000000000";
--ram(86) <= "00000000101000110011000000010010";
--ram(87) <= "00000000101000110011100000010100";
--ram(88) <= "00000000111001100011100000010100";
--ram(89) <= "00100000000001110000000000110000";
--ram(90) <= "00100000000001010000000000110001";
--ram(91) <= "00011100000010100000000000101111";
--ram(92) <= "00011100000010110000000000110000";
--ram(93) <= "00011100000011000000000000110001";
--ram(94) <= "00000001010011000110100000010010";
--ram(95) <= "00101000000011010000000000001001";
--ram(96) <= "00001001101011100000000000100000";
--ram(97) <= "00011100000011110000000000110000";
--ram(98) <= "00010101011010110000000000000001";
--ram(99) <= "00001001101011010000000000000001";
--ram(100) <= "00101100000011011111111111111101";
--ram(101) <= "00011001111011110000000000000001";
--ram(102) <= "00000101110011100000000000000001";
--ram(103) <= "00101100000011101111111111111101";
--ram(104) <= "00000001111010110101100000010011";
--ram(105) <= "00000001000010000100000000010000";
--ram(106) <= "00011101000010010000000000001110";
--ram(107) <= "00000001001010110001100000010000";
--ram(108) <= "00000100011000110000000000000000";
--ram(109) <= "00000000101000110011000000010010";
--ram(110) <= "00000000101000110011100000010100";
--ram(111) <= "00000000111001100011100000010100";
--ram(112) <= "00100000000001110000000000110000";
--ram(113) <= "00100000000000110000000000110001";
--ram(114) <= "00011100000010100000000000101111";
--ram(115) <= "00011100000010110000000000110000";
--ram(116) <= "00011100000011000000000000110001";
--ram(117) <= "00000001010011000110100000010010";
--ram(118) <= "00101000000011010000000000001001";
--ram(119) <= "00001001101011100000000000100000";
--ram(120) <= "00011100000011110000000000110000";
--ram(121) <= "00010101011010110000000000000001";
--ram(122) <= "00001001101011010000000000000001";
--ram(123) <= "00101100000011011111111111111101";
--ram(124) <= "00011001111011110000000000000001";
--ram(125) <= "00000101110011100000000000000001";
--ram(126) <= "00101100000011101111111111111101";
--ram(127) <= "00000001111010110101100000010011";
--ram(128) <= "00000101000010000000000000000001";
--ram(129) <= "00011101000010010000000000001110";
--ram(130) <= "00000001001010110010100000010000";
--ram(131) <= "00000100101001010000000000000000";
--ram(132) <= "00000100001000010000000000000001";
--ram(133) <= "00101110100000011111111111010010";
--ram(134) <= "00000100000000010000000000000000";
--ram(135) <= "00100000001000110000000000101101";
--ram(136) <= "00000100011000110000000000000000";
--ram(137) <= "00000100001000010000000000000001";
--ram(138) <= "00100000001001010000000000101101";
--ram(139) <= "00000100101001010000000000000000";
--ram(140) <= "00000100000000010000000000000000";
--ram(141) <= "00011100001000110000000000101101";
--ram(142) <= "00000100001000010000000000000001";
--ram(143) <= "00011100001001010000000000101101";
--ram(144) <= "00000100000100000000000000000001";
--ram(145) <= "00000100000000010000000000001100";
--ram(146) <= "00000100001000100000000000000000";
--ram(147) <= "00000000001000010000100000010000";
--ram(148) <= "00000100001000010000000000000001";
--ram(149) <= "00011100001001100000000000001110";
--ram(150) <= "00000000110001010010100000010001";
--ram(151) <= "00100000000001010000000000110000";
--ram(152) <= "00100000000000110000000000110001";
--ram(153) <= "00011100000010100000000000101111";
--ram(154) <= "00011100000010110000000000110000";
--ram(155) <= "00011100000011000000000000110001";
--ram(156) <= "00000001010011000110100000010010";
--ram(157) <= "00101000000011010000000000001001";
--ram(158) <= "00001001101011100000000000100000";
--ram(159) <= "00011100000011110000000000110000";
--ram(160) <= "00011001011010110000000000000001";
--ram(161) <= "00001001101011010000000000000001";
--ram(162) <= "00101100000011011111111111111101";
--ram(163) <= "00010101111011110000000000000001";
--ram(164) <= "00000101110011100000000000000001";
--ram(165) <= "00101100000011101111111111111101";
--ram(166) <= "00000001111010110101100000010011";
--ram(167) <= "00000000011010110100000000010010";
--ram(168) <= "00000000011010110011100000010100";
--ram(169) <= "00000000111010000010100000010100";
--ram(170) <= "00001000001000010000000000000001";
--ram(171) <= "00011100001001100000000000001110";
--ram(172) <= "00000000110000110001100000010001";
--ram(173) <= "00100000000000110000000000110000";
--ram(174) <= "00100000000001010000000000110001";
--ram(175) <= "00011100000010100000000000101111";
--ram(176) <= "00011100000010110000000000110000";
--ram(177) <= "00011100000011000000000000110001";
--ram(178) <= "00000001010011000110100000010010";
--ram(179) <= "00101000000011010000000000001001";
--ram(180) <= "00001001101011100000000000100000";
--ram(181) <= "00011100000011110000000000110000";
--ram(182) <= "00011001011010110000000000000001";
--ram(183) <= "00001001101011010000000000000001";
--ram(184) <= "00101100000011011111111111111101";
--ram(185) <= "00010101111011110000000000000001";
--ram(186) <= "00000101110011100000000000000001";
--ram(187) <= "00101100000011101111111111111101";
--ram(188) <= "00000001111010110101100000010011";
--ram(189) <= "00000000101010110100000000010010";
--ram(190) <= "00000000101010110011100000010100";
--ram(191) <= "00000000111010000001100000010100";
--ram(192) <= "00001000001000010000000000000001";
--ram(193) <= "00101110000000011111111111010010";
--ram(194) <= "00011100001001100000000000001110";
--ram(195) <= "00000000110001010010100000010001";
--ram(196) <= "00001000001000010000000000000001";
--ram(197) <= "00011100001001100000000000001110";
--ram(198) <= "00000000110000110001100000010001";
--ram(199) <= "00100000000000110000000000101011";
--ram(200) <= "00000100011000110000000000000000";
--ram(201) <= "00100000000001010000000000101100";
--ram(202) <= "00000100101001010000000000000000";
--
--
----			ram(0) <= "00000100000000010000000000000111";
----			ram(1) <= "00000100000000100000000000001000";
----			ram(2) <= "00000000010000010001100000010000";
----			ram(0) <= "00100100000000010000000000000100"; -- beq
----			ram(0) <= "00101000000000010000000000000010"; -- load
----			ram(1) <= "00000100001001000000000000000000"; -- addi
----			ram(1) <= "00000100000000010000000000000010";
----			ram(2) <= "00000100000000110000000000001010";
----			ram(3) <= "00000100000001000000000000001110";
----			ram(4) <= "00000100000001010000000000000010";
----			ram(5) <= "00100000011001000000000000000010";
----			ram(6) <= "00100000011000110000000000000001";
----			ram(7) <= "00000000011001000010000000010001";
----			ram(8) <= "00001000000001000000000000000001";
----			ram(9) <= "00000000011000100010000000010010";
----			ram(10) <= "00001100010001000000000000001010";
----			ram(11) <= "00000000011000100010000000010011";
----			ram(12) <= "00011100011000100000000000000001";
----			ram(13) <= "00010000010001000000000000001010";
----			ram(14) <= "00000000011000100010000000010100";
----			ram(15) <= "00010100010001000000000000001010";
----			ram(16) <= "00011000010001000000000000001010";
----			ram(17) <= "00101000000001011111111111111110";
----			ram(18) <= "00100100100001010000000000000000";
----			ram(19) <= "00101100100001010000000000000000";
----			ram(20) <= "00110000000000000000000000010101";
----			ram(21) <= "11111100000000000000000000000000";

 		END IF;
	END PROCESS;
	
	instr <= ram(CONV_INTEGER(read_addr));	

	
end Behavioral;

